/**
 * PyObjectWrapper.svh
 *
 * Copyright 2024 Matthew Ballance and Contributors
 *
 * Licensed under the Apache License, Version 2.0 (the "License"); you may 
 * not use this file except in compliance with the License.  
 * You may obtain a copy of the License at:
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software 
 * distributed under the License is distributed on an "AS IS" BASIS, 
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  
 * See the License for the specific language governing permissions and 
 * limitations under the License.
 *
 * Created on:
 *     Author: 
 */
class PyObjectWrapper;
    PyObject            m_hndl;
    bit                 m_owned;

    function new(PyObject hndl, bit owned=1);
        m_hndl = hndl;
    endfunction

    function longint unsigned getAttrUi64(string name);
    endfunction

    function void setAttrUi64(string name, longint unsigned val);
    endfunction

//    static function PyObjectWrapper newClass()

endclass

