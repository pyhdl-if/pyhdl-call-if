
module smoke;

  initial begin
    $display("smoke");
  end
endmodule
